`include "lisnoc_def.vh"

`undef FLIT_WIDTH

`undef FLIT_TYPE_MSB
`undef FLIT_TYPE_WIDTH
`undef FLIT_TYPE_LSB

`undef FLIT_CONTENT_WIDTH
`undef FLIT_CONTENT_MSB
`undef FLIT_CONTENT_LSB

`undef FLIT_DEST_WIDTH
`undef FLIT_DEST_MSB
`undef FLIT_DEST_LSB

`undef PACKET_CLASS_MSB
`undef PACKET_CLASS_WIDTH
`undef PACKET_CLASS_LSB

`undef PACKET_CLASS_DMA

// source address field  of header flit
`undef SOURCE_MSB
`undef SOURCE_WIDTH
`undef SOURCE_LSB

// packet id field  of header flit
`undef PACKET_ID_MSB  
`undef PACKET_ID_WIDTH 
`undef PACKET_ID_LSB  

`undef PACKET_TYPE_MSB   
`undef PACKET_TYPE_WIDTH 
`undef PACKET_TYPE_LSB   

`undef PACKET_TYPE_L2R_REQ 
`undef PACKET_TYPE_R2L_REQ 
`undef PACKET_TYPE_L2R_RESP
`undef PACKET_TYPE_R2L_RESP

`undef PACKET_REQ_LAST
`undef PACKET_RESP_LAST

`undef SIZE_MSB   
`undef SIZE_WIDTH 
`undef SIZE_LSB  

`undef DMA_REQUEST_WIDTH 

`undef DMA_REQFIELD_LADDR_WIDTH
`undef DMA_REQFIELD_SIZE_WIDTH
`undef DMA_REQFIELD_RTILE_WIDTH
`undef DMA_REQFIELD_RADDR_WIDTH

`undef DMA_REQFIELD_LADDR_MSB 
`undef DMA_REQFIELD_LADDR_LSB 
`undef DMA_REQFIELD_SIZE_MSB  
`undef DMA_REQFIELD_SIZE_LSB  
`undef DMA_REQFIELD_RTILE_MSB 
`undef DMA_REQFIELD_RTILE_LSB 
`undef DMA_REQFIELD_RADDR_MSB 
`undef DMA_REQFIELD_RADDR_LSB 
`undef DMA_REQFIELD_DIR       

`undef DMA_REQUEST_INVALID 
`undef DMA_REQUEST_VALID   

`undef DMA_REQMASK_WIDTH 
`undef DMA_REQMASK_LADDR 
`undef DMA_REQMASK_SIZE  
`undef DMA_REQMASK_RTILE 
`undef DMA_REQMASK_RADDR 
`undef DMA_REQMASK_DIR   
