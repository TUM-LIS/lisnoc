/**
 * This file is part of LISNoC.
 * 
 * LISNoC is free hardware: you can redistribute it and/or modify
 * it under the terms of the GNU Lesser General Public License as 
 * published by the Free Software Foundation, either version 3 of 
 * the License, or (at your option) any later version.
 *
 * As the LGPL in general applies to software, the meaning of
 * "linking" is defined as using the LISNoC in your projects at
 * the external interfaces.
 * 
 * LISNoC is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU Lesser General Public 
 * License along with LISNoC. If not, see <http://www.gnu.org/licenses/>.
 * 
 * =================================================================
 * 
 * This file should be included at the end of every file that
 * includes lisnoc_def.vh. It avoids any conflicts with your system.
 *
 * (c) 2011-2012 by the author(s)
 * 
 * Author(s): 
 *    Stefan Wallentowitz, stefan.wallentowitz@tum.de
 *    Andreas Lankes, andreas.lankes@tum.de
 *    Michael Tempelmeier, michael.tempelmeier@tum.de
 */

`undef FLIT_TYPE_PAYLOAD
`undef FLIT_TYPE_HEADER
`undef FLIT_TYPE_LAST
`undef FLIT_TYPE_SINGLE

`undef SELECT_NORTH
`undef SELECT_EAST
`undef SELECT_SOUTH
`undef SELECT_WEST
`undef SELECT_LOCAL

`undef NORTH
`undef EAST
`undef SOUTH
`undef WEST
`undef LOCAL

